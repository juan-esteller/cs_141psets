----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    12:02:52 09/16/2017 
-- Design Name: 
-- Module Name:    mux_16to1 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity mux_16to1 is
    Port ( I_0 : in  STD_LOGIC;
           I_1 : in  STD_LOGIC;
           I_2 : in  STD_LOGIC;
           I_3 : in  STD_LOGIC;
           I_4 : in  STD_LOGIC;
           I_5 : in  STD_LOGIC;
           I_6 : in  STD_LOGIC;
           I_7 : in  STD_LOGIC;
           I_8 : in  STD_LOGIC;
           I_9 : in  STD_LOGIC;
           I_10 : in  STD_LOGIC;
           I_11 : in  STD_LOGIC;
           I_12 : in  STD_LOGIC;
           I_13 : in  STD_LOGIC;
           I_14 : in  STD_LOGIC;
           I_15 : in  STD_LOGIC;
           control : in  STD_LOGIC;
           result : out  STD_LOGIC);
end mux_16to1;

architecture Behavioral of mux_16to1 is

begin


end Behavioral;

